-------------------------------------------------------------------------------
-- Title      : twominus scan logic
-- Project    : 
-------------------------------------------------------------------------------
-- File       : twominus_scan.vhd
-- Author     : sdong  <sdong@sdong-ubuntu>
-- Company    : 
-- Created    : 2021-10-21
-- Last update: 2021-10-21
-- Platform   : 
-- Standard   : VHDL'2008
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2021 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-10-21  1.0      sdong   Created
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity twominus_scan is
  port (
    clk : in std_logic;  -- The twominus clock is generated by one MMMC, and the frequency is controlled by the software.
    rst : in std_logic;

    start_scan : in  std_logic;         -- Start signal from software
    reset_scan : in  std_logic;
    -- The io ports of the ASIC
    speak      : out std_logic;
    start      : out std_logic;
    rst_out    : out std_logic
    );
end twominus_scan;

architecture behv of twominus_scan is
  -- declarative_items (signal declarations, component declarations, etc.)  
  type SCAN_STATE is (IDLE, RESET_CHIP, ASS_START, ASS_SPEAK);
  signal state_reg, state_next : SCAN_STATE;

  signal rst_cnt : integer range 0 to 3;

  --Debug
  attribute mark_debug               : string;
  attribute mark_debug of rst_cnt    : signal is "true";
  attribute mark_debug of speak      : signal is "true";
  attribute mark_debug of start      : signal is "true";
  attribute mark_debug of rst_out    : signal is "true";
  attribute mark_debug of start_scan : signal is "true";
  attribute mark_debug of reset_scan : signal is "true";

begin
  -- architecture body

  process(clk, rst)
  begin
    if rst = '1' then
      state_reg <= IDLE;
    elsif rising_edge(clk) then
      state_reg <= state_next;
    end if;
  end process;

  process(all)
  begin
    state_next <= state_reg;
    case state_reg is
      when IDLE =>
        if ?? start_scan then
          state_next <= RESET_CHIP;
        end if;
      when RESET_CHIP =>
        if rst_cnt = 3 then
          state_next <= ASS_START;
        end if;
      when ASS_START =>
        state_next <= ASS_SPEAK;
      when ASS_SPEAK =>
        if ?? reset_scan then
          state_next <= IDLE;
        end if;
      when others =>
        state_next <= IDLE;
    end case;
  end process;

  process(clk)
  begin
    if rising_edge(clk) then
      case(state_next) is
        when IDLE =>
          speak   <= '0';
          start   <= '0';
          rst_out <= '0';
          rst_cnt <= 0;
        when RESET_CHIP =>
          rst_out <= '1';
          rst_cnt <= rst_cnt + 1;
        when ASS_START =>
          rst_out <= '0';
          start   <= '1';
          rst_cnt <= 0;
        when ASS_SPEAK =>
          start   <= '0';
          speak   <= '1';
          rst_cnt <= 0;
        when others => null;
      end case;
    end if;
  end process;

end behv;
